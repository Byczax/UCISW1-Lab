----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:17:17 12/01/2021 
-- Design Name: 
-- Module Name:    gfunctiontruthtable - Dataflow 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity gfunctiontruthtable is
    Port ( WEJ : in  STD_LOGIC_VECTOR (3 downto 0);
           WYJ : out  STD_LOGIC);
end gfunctiontruthtable;

architecture Dataflow of gfunctiontruthtable is

begin
	with WEJ select
	WYJ <= '1' when "0001" | "0101" | "1000" | "1010" | "1110",
			 '0' when others;

end Dataflow;

